module andgate (c,a,b);
input a,b;
output c;
and a1(c,a,b);  

endmodule

